package bloom_filter_regs_pkg;

// Registers:
parameter EN             = 0;
parameter HASH_LUT_CLEAN = 1;
parameter BASIC_REGS_CNT = 2;

endpackage
